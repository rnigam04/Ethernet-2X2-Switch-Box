//This conist of the SV testbench for Ethernet 2X2 Switch Box
// All the details were present in the README File
module ethernetswbox_tb();

endmodule // ethernetswbox_tb
